//============================================================================//
//    FCUDA
//    Copyright (c) <2016> 
//    <University of Illinois at Urbana-Champaign>
//    <University of California at Los Angeles> 
//    All rights reserved.
// 
//    Developed by:
// 
//        <ES CAD Group & IMPACT Research Group>
//            <University of Illinois at Urbana-Champaign>
//            <http://dchen.ece.illinois.edu/>
//            <http://impact.crhc.illinois.edu/>
// 
//        <VAST Laboratory>
//            <University of California at Los Angeles>
//            <http://vast.cs.ucla.edu/>
// 
//        <Hardware Research Group>
//            <Advanced Digital Sciences Center>
//            <http://adsc.illinois.edu/>
//============================================================================//

`timescale 1ns / 1ps
`include "noc_pkt.vh" 

// The module implementing the directory
// There are two implementations: one uses not-real many-ported BRAMs, the
// other uses a single BRAM that has arbitration for ports
module dirnew(

  input wire clk,
  input wire rst,

  input  wire [`DIR_READEN_WIDTH      - 1: 0] readen,
  input  wire [`TOTAL_TAG_WIDTH       - 1: 0] tags,
  input  wire [`TOTAL_INDEX_WIDTH     - 1: 0] indecies,
  input  wire [`TOTAL_ROUTER_ID_WIDTH - 1: 0] router_ids,
  input  wire [`TOTAL_PKT_TYPE_WIDTH  - 1: 0] pkt_types,
  input  wire [`TOTAL_SRC_ADDR_WIDTH  - 1: 0] src_addrs,
  `ifdef ENABLE_OUTSTANDING_ARRAY
  input  wire [`TOTAL_DEST_ADDR_WIDTH  - 1: 0] dest_addrs,
  input  wire [`NUM_INPUTS - 1 : 0] wasreplaced,
`endif
input  wire [`NUM_INPUTS - 1 : 0] pkt_valids,
output wire [`DIR_READEN_WIDTH      - 1: 0] hits,
output wire [`TOTAL_RESULT_SIZE     - 1: 0] results
);

parameter [`ROUTER_ID_WIDTH-1:0] ROUTER_ID = {`ROUTER_ID_WIDTH{1'b0}};

`ifdef REAL_DIRECTORY_IMPLEMENTATION   // New directory implementation that uses arbitration on a real 2-ported BRAM

// contents of single directory entry == tag + dest + valid
localparam BRAM_SIZE = `TAG_WIDTH + `DESTWIDTH + 1;

// BRAM writeenable
wire we1;
wire we2;

// BRAM index
wire [`INDEX_WIDTH-1:0] addr1;
wire [`INDEX_WIDTH-1:0] addr2;

// BRAM input
wire [BRAM_SIZE-1:0] di1;
wire [BRAM_SIZE-1:0] di2;

// BRAM output
wire [BRAM_SIZE-1:0] do1;
wire [BRAM_SIZE-1:0] do2;

// choose which input port to allow to read/write directory
wire [1 : 0]  sel1;
wire sel2;

// this BRAM contains the directory
bram #(
  .DATASIZE(BRAM_SIZE),
  .ADDRWIDTH(`INDEX_WIDTH),
  .DEPTH(`DIRECTORY_SIZE)
) dbram (  
  .clk(clk),    // done
  .rst(rst),    // done
  .we1(we1),     // done
  .we2(we2),     // done
  .addr1(addr1), // done
  .addr2(addr2), // done
  .di1(di1),     // done
  .di2(di2),     // done
  .do1(do1),     // done
  .do2(do2)      // done
);


//   {x,y,x}0 ==> readenable for input port 0,1,2 (x,y,z)
//   {x,y,x}1 ==> writeenable for input port 0,1,2 (x,y,z)  
wire X0, X1;
wire Y0, Y1; 
wire Z0, Z1;

// bits 1,0 of counter
wire C1, C0;

// output: generates select bits to choose which port gets access
wire S1, S0; 

// In arbitration scheme, writes to directory have priority over reads. This
// can be experimented with. 

// arbitration is done by round-robin counters
reg [1:0] ctr1;  // counts 0,1,2,0,1,2,...
reg ctr2;        // counts 0,1,0,1,0,1,...

assign X0 = readen[0];
assign X1 = check_we (0, router_ids, pkt_types,pkt_valids); 
assign Y0 = readen[1];
assign Y1 = check_we (1, router_ids, pkt_types,pkt_valids); 
assign Z0 = readen[2];
assign Z1 = check_we (2, router_ids, pkt_types,pkt_valids); 

assign C0 = ctr1[1];
assign C1 = ctr1[0];


// arbitration counters
always @(posedge clk)
begin
  if (rst) begin
    ctr1 <= 0;
    ctr2 <= 0;
  end else begin
    if (ctr1 == 2) begin
      ctr1 <= 0;
    end else begin
      ctr1 <= ctr1 + 1;
    end
    ctr2 <= ctr2 + 1;
  end
end

// logic generated by bont scripts
assign S1=Z1&(!Z0)&C1&(!C0) |X0&Z1&(!Z0)&(!C0) |(!X1)&Z1&(!Z0)&(!C0) |X0&Y0&Z1&(!Z0)&(!C1) |(!X1)&Y0&Z1&(!Z0)&(!C1) |X0&(!Y1)&Z1&(!Z0)&(!C1) |(!X1)&(!Y1)&Z1&(!Z0)&(!C1) |X0&Y0&(!Z1)&Z0&C1&(!C0) |X1&X0&(!Y1)&(!Z1)&Z0&(!C0) |(!X1)&(!Y1)&(!Z1)&Z0&C1&(!C0) |(!X1)&(!X0)&Y0&(!Z1)&Z0&(!C0) |X1&X0&Y1&Y0&(!Z1)&Z0&(!C1) |(!X1)&(!X0)&Y1&Y0&(!Z1)&Z0&(!C1) |X1&X0&(!Y1)&(!Y0)&(!Z1)&Z0&(!C1) |(!X1)&(!X0)&(!Y1)&(!Y0)&(!Z1)&Z0&(!C1);

assign S0=Y1&(!Y0)&(!C1)&C0 |X0&Y1&(!Y0)&Z0&(!C0) |(!X1)&Y1&(!Y0)&Z0&(!C0) |X0&Y1&(!Y0)&(!Z1)&(!C0) |(!X1)&Y1&(!Y0)&(!Z1)&(!C0) |X0&(!Y1)&Y0&Z0&(!C1)&C0 |(!X1)&(!Y1)&Y0&Z0&(!C1)&C0 |X0&(!Y1)&Y0&(!Z1)&(!C1)&C0 |(!X1)&(!Y1)&Y0&(!Z1)&(!C1)&C0 |X1&X0&(!Y1)&Y0&Z1&Z0&(!C0) |(!X1)&(!X0)&(!Y1)&Y0&Z1&Z0&(!C0) |X1&X0&(!Y1)&Y0&(!Z1)&(!Z0)&(!C0) |(!X1)&(!X0)&(!Y1)&Y0&(!Z1)&(!Z0)&(!C0);

wire A0,A1,B0,B1,C;

// readen and we for ports 3, 4
assign A0 = readen[3]; 
assign A1 = check_we (3, router_ids, pkt_types,pkt_valids); 
assign B0 = readen[4];
assign B1 = check_we (4, router_ids, pkt_types,pkt_valids); 

// short name for counter value -
assign C = ctr2;

// result bit -- choose [4] or [5]
wire S;

assign S=B1&(!B0)&C |A0&B1&(!B0) |(!A1)&B1&(!B0) |A0&(!B1)&B0&C |A1&A0&(!B1)&B0 |(!A1)&(!A0)&(!B1)&B0;


// assign select bits based on output of above logic
// this logic is pretty expensive...
//   Or not -- e.g. LUTs have 6 inputs and can implement any function => maybe
//   only 1 lut?
assign sel1[1] = S1;
assign sel1[0] = S0;
assign sel2 = S;

// all that is left is to assign sel1, sel2
// do this based on output of the combinational logic
reg [1:0] sel1_reg;
reg sel2_reg;

reg[`DIR_READEN_WIDTH      - 1: 0]  readen_reg;
reg[`TOTAL_TAG_WIDTH       - 1: 0]  tags_reg;

always @(posedge clk) 
begin
  sel1_reg <= sel1;
  sel2_reg <= sel2;
  readen_reg <= readen;
  tags_reg <= tags;
end

`ifdef ENABLE_OUTSTANDING_ARRAY
reg[`NUM_INPUTS-1:              0]  wasreplaced_reg;
reg[`TOTAL_DEST_ADDR_WIDTH  - 1: 0] dest_addrs_reg;
always @(posedge clk) 
begin
  dest_addrs_reg  <= dest_addrs;
  wasreplaced_reg <= wasreplaced;
end
`endif // ENABLE_OUTSTANDING_ARRAY

genvar k;

// the following assigns output results per-port based on tag match, valid,
// and whether or not given input was selected and was being read
// FIXME: changed to remove reg delay...this seems so wrong, though...
`ifdef ENABLE_OUTSTANDING_ARRAY
generate 
  for (k =0; k < 3; k = k + 1) begin:RESULTS1
    // 
    assign hits[k] = ((sel1_reg== k) & (do1[BRAM_SIZE-1]) & (readen_reg[k] == 1'b1) & 
    (tags_reg[`BOUNDS(k,`TAG_WIDTH)] == do1[`DESTWIDTH + `TAG_WIDTH -1 : `DESTWIDTH])) | 
    wasreplaced_reg[k];

    assign results[`BOUNDS(k,`DESTWIDTH)] = wasreplaced_reg[k] ? dest_addrs_reg[`BOUNDS(k,`DESTWIDTH)] : do1[`DESTWIDTH-1:0];
  end

  for (k =3; k < `NUM_INPUTS; k = k + 1) begin:RESULTS2
    assign hits[k] = ((sel2_reg== (k - 3)) & (do2[BRAM_SIZE-1])  & (readen_reg[k] == 1'b1) & 
    (tags_reg[`BOUNDS(k,`TAG_WIDTH)] == do2[`DESTWIDTH + `TAG_WIDTH -1 : `DESTWIDTH])) |
    wasreplaced_reg[k];

    assign results[`BOUNDS(k,`DESTWIDTH)] = wasreplaced_reg[k] ? dest_addrs_reg[`BOUNDS(k,`DESTWIDTH)] : do2[`DESTWIDTH-1:0];
  end
endgenerate
`else
generate 
  for (k =0; k < 3; k = k + 1) begin:RESULTS1
    assign hits[k] = ((sel1_reg== k) & (do1[BRAM_SIZE-1]) & (readen_reg[k] == 1'b1) & 
    (tags_reg[`BOUNDS(k,`TAG_WIDTH)] == do1[`DESTWIDTH + `TAG_WIDTH -1 : `DESTWIDTH]));

    assign results[`BOUNDS(k,`DESTWIDTH)] = do1[`DESTWIDTH-1:0];
  end

  for (k =3; k < `NUM_INPUTS; k = k + 1) begin:RESULTS2
    assign hits[k] = ((sel2_reg== (k - 3)) & (do2[BRAM_SIZE-1])  & (readen_reg[k] == 1'b1) & 
    (tags_reg[`BOUNDS(k,`TAG_WIDTH)] == do2[`DESTWIDTH + `TAG_WIDTH -1 : `DESTWIDTH]));

    assign results[`BOUNDS(k,`DESTWIDTH)] = do2[`DESTWIDTH-1:0];
  end
endgenerate
`endif


// (ROUTER_ID == router_ids[`BOUNDS(0,`ROUTER_ID_WIDTH)] && `TYPE_RESPONSE_ADDR ==  pkt_types [`BOUNDS(0,`DATA_TYPEWIDTH)])

// set writeenable for BRAM port 0

// assign we1 = (sel1 == 2'b00) ? check_we(0, router_ids, pkt_types) :
//              (sel1 == 2'b01) ? check_we(1, router_ids, pkt_types) : 
//              (sel1 == 2'b10) ? check_we(2, router_ids, pkt_types) :  0; // 0 if (sel = 11)

assign we1 = (sel1 == 2'b00) ? X1 :
(sel1 == 2'b01) ? Y1 : 
(sel1 == 2'b10) ? Z1 :  0; // 0 if (sel = 11)

// set writeenable for BRAM port 1
// assign we2 = (sel2 == 1'b0) ? check_we(3,router_ids, pkt_types) :
//              (sel2 == 1'b1) ? check_we(4,router_ids, pkt_types) :     0; // 0 if (sel == ??)

assign we2 = (sel2 == 1'b0) ? A1 :
(sel2 == 1'b1) ? B1 :     0; // 0 if (sel == ??)


// assign di1 as { valid, tag, data}
assign di1 = (sel1 == 2'b00) ? {1'b1, tags[`BOUNDS(0,`TAG_WIDTH)], src_addrs[`BOUNDS(0,`DATA_SRCWIDTH)] }:
(sel1 == 2'b01) ? {1'b1, tags[`BOUNDS(1,`TAG_WIDTH)], src_addrs[`BOUNDS(1,`DATA_SRCWIDTH)] }: 
(sel1 == 2'b10) ? {1'b1, tags[`BOUNDS(2,`TAG_WIDTH)], src_addrs[`BOUNDS(2,`DATA_SRCWIDTH)] }:  0; // 0 if (sel = 11)

// assign di1 as { valid, tag, data}
assign di2 = (sel2 == 1'b0) ? {1'b1, tags[`BOUNDS(3,`TAG_WIDTH)], src_addrs[`BOUNDS(3,`DATA_SRCWIDTH)] }:
(sel2 == 1'b1) ? {1'b1, tags[`BOUNDS(4,`TAG_WIDTH)], src_addrs[`BOUNDS(4,`DATA_SRCWIDTH)] }:     0; // 0 if (sel == ??)

// choose BRAM index for port 0
assign addr1 = (sel1 == 2'b00) ? indecies  [`BOUNDS(0,`INDEX_WIDTH)]:
(sel1 == 2'b01) ? indecies  [`BOUNDS(1,`INDEX_WIDTH)]: 
(sel1 == 2'b10) ? indecies  [`BOUNDS(2,`INDEX_WIDTH)]:  0; // 0 if (sel = 11)

// choose BRAM index for port 1
assign addr2 = (sel2 == 1'b0) ? indecies  [`BOUNDS(3,`INDEX_WIDTH)]:
(sel2 == 1'b1) ? indecies  [`BOUNDS(4,`INDEX_WIDTH)]:     0; // 0 if (sel == ??)

function check_we;
    input [31:0] input_id;
    input  [`TOTAL_ROUTER_ID_WIDTH - 1: 0] router_ids;
    input  [`TOTAL_PKT_TYPE_WIDTH  - 1: 0] pkt_types;
    input  [`NUM_INPUTS  - 1: 0] pkt_valids;
  begin
    check_we = (pkt_valids[input_id]) & ((ROUTER_ID == router_ids[(input_id + 1) * `ROUTER_ID_WIDTH -1 -: `ROUTER_ID_WIDTH]) & (`TYPE_RESPONSE_ADDR ==  pkt_types [(input_id + 1)*`DATA_TYPEWIDTH -1 -: `DATA_TYPEWIDTH]));
  end
endfunction

`else // Original many-ported directory implementation

// caches
reg [`DESTWIDTH-1:0]      data_array [`DIRECTORY_SIZE-1:0];
reg [`TAG_WIDTH-1:0]      tag_array  [`DIRECTORY_SIZE-1:0];
reg [`DIRECTORY_SIZE-1:0] valid_array  ; /* just one bit */

// .......
wire [`INDEX_WIDTH-1:0]   cur_index_arr [`NUM_INPUTS-1:0]  ;
wire [`DATA_SRCWIDTH-1:0] cur_data_arr [`NUM_INPUTS-1:0]  ;
wire [`TAG_WIDTH-1:0]     cur_tag_arr [`NUM_INPUTS-1:0]  ;

wire wr_en[`NUM_INPUTS-1:0];

/* initializes valid bits to 0 */
integer arrayinit;
initial begin
  for(arrayinit=0;arrayinit<`DIRECTORY_SIZE;arrayinit = arrayinit + 1) begin
    valid_array[arrayinit] = 1'b0;
  end
end

integer j;

integer num_cache_insertions;

always @(posedge clk or posedge rst) begin
  if (rst) begin
    num_cache_insertions = 0;
  end else begin
    for (j = 0; j < `NUM_INPUTS; j = j + 1) begin
      if (wr_en[j] == 1'b1) begin
        num_cache_insertions = num_cache_insertions + 1;
        tag_array[cur_index_arr[j]]   = cur_tag_arr[j];
        data_array[cur_index_arr[j]]  = cur_data_arr[j];
        valid_array[cur_index_arr[j]] = 1'b1;
      end
    end
  end
end

genvar i;
generate
  for (i =0; i < `NUM_INPUTS; i = i + 1) begin:ARRAYACCESS
    wire [`TAG_WIDTH-1:0]         cur_tag;
    wire [`ROUTER_ID_WIDTH-1:0]   cur_router_id;
    wire [`INDEX_WIDTH-1:0]       cur_index;
    wire [`DATA_TYPEWIDTH-1:0]    cur_type;
    wire [`DATA_SRCWIDTH-1:0]     cur_src_addr;

    wire [`TAG_WIDTH-1:0]   match_tag; 

    // rip off bits from input
    assign cur_router_id = router_ids[`BOUNDS(i,`ROUTER_ID_WIDTH)];
    assign cur_tag       = tags      [`BOUNDS(i,`TAG_WIDTH)];
    assign cur_index     = indecies  [`BOUNDS(i,`INDEX_WIDTH)];
    assign cur_type      = pkt_types [`BOUNDS(i,`DATA_TYPEWIDTH)];
    assign cur_src_addr  = src_addrs [`BOUNDS(i,`DATA_SRCWIDTH)];



    `ifdef ENABLE_OUTSTANDING_ARRAY
    wire [`DESTWIDTH-1:0]         cur_dest_addr;
    assign cur_dest_addr = dest_addrs[`BOUNDS(i,`DESTWIDTH)];
    `endif

    // decide to write cache or not
    assign wr_en[i]         = cur_router_id == ROUTER_ID && cur_type == `TYPE_RESPONSE_ADDR;

    // set bits for cache lookup (or write)
    assign cur_index_arr[i] = cur_index;
    assign cur_tag_arr[i]   = cur_tag;
    assign cur_data_arr[i]  = cur_src_addr;

    // lookup in tag array
    assign match_tag = tag_array[cur_index];

    // check for hit
    `ifdef ENABLE_OUTSTANDING_ARRAY
    assign hits[i] = ((cur_tag == match_tag) & valid_array[cur_index] & readen[i]) | wasreplaced[i];
    assign results[`BOUNDS(i,`DESTWIDTH)] = wasreplaced[i] ? cur_dest_addr  : data_array[cur_index];
    `else
    assign hits[i] = ((cur_tag == match_tag) & valid_array[cur_index] & readen[i]);
    assign results[`BOUNDS(i,`DESTWIDTH)] = data_array[cur_index];
    `endif
  end
endgenerate
`endif

endmodule
